module registerFile
(
  input [4:0] RS1,
  input [4:0] RS2,
  input [4:0] RD,
  input [63:0] WriteData,
  output reg [63:0] ReadData1,
  output reg [63:0] ReadData2,
  input clk, reset, RegWrite
);

  reg [63:0] Registers [31:0];
  
  initial
  begin
  Registers[0] <= 64'b00000000000000000000000000000000000000000000000000000000000000;
  Registers[1] <= 64'b00000000000000000000000000000000000000000000000000000000000001;
  Registers[2] <= 64'b00000000000000000000000000000000000000000000000000000000000010;
  Registers[3] <= 64'b00000000000000000000000000000000000000000000000000000000000011;
  Registers[4] <= 64'b00000000000000000000000000000000000000000000000000000000000100;
  Registers[5] <= 64'b00000000000000000000000000000000000000000000000000000000000101;
  Registers[6] <= 64'b00000000000000000000000000000000000000000000000000000000000110;
  Registers[7] <= 64'b00000000000000000000000000000000000000000000000000000000000111;
  Registers[8] <= 64'b00000000000000000000000000000000000000000000000000000000001000;
  Registers[9] <= 64'b00000000000000000000000000000000000000000000000000000000001001;
  Registers[10] <= 64'b00000000000000000000000000000000000000000000000000000000001010;
  Registers[11] <= 64'b00000000000000000000000000000000000000000000000000000000001011;
  Registers[12] <= 64'b00000000000000000000000000000000000000000000000000000000001100;
  Registers[13] <= 64'b00000000000000000000000000000000000000000000000000000000001101;
  Registers[14] <= 64'b00000000000000000000000000000000000000000000000000000000001110;
  Registers[15] <= 64'b00000000000000000000000000000000000000000000000000000000001111;
  Registers[16] <= 64'b00000000000000000000000000000000000000000000000000000000010000;
  Registers[17] <= 64'b00000000000000000000000000000000000000000000000000000000010001;
  Registers[18] <= 64'b00000000000000000000000000000000000000000000000000000000010010;
  Registers[19] <= 64'b00000000000000000000000000000000000000000000000000000000010011;
  Registers[20] <= 64'b00000000000000000000000000000000000000000000000000000000010100;
  Registers[21] <= 64'b00000000000000000000000000000000000000000000000000000000010101;
  Registers[22] <= 64'b00000000000000000000000000000000000000000000000000000000010110;
  Registers[23] <= 64'b00000000000000000000000000000000000000000000000000000000010111;
  Registers[24] <= 64'b00000000000000000000000000000000000000000000000000000000011000;
  Registers[25] <= 64'b00000000000000000000000000000000000000000000000000000000011001;
  Registers[26] <= 64'b00000000000000000000000000000000000000000000000000000000011010;
  Registers[27] <= 64'b00000000000000000000000000000000000000000000000000000000011011;
  Registers[28] <= 64'b00000000000000000000000000000000000000000000000000000000011100;
  Registers[29] <= 64'b00000000000000000000000000000000000000000000000000000000011101;
  Registers[30] <= 64'b00000000000000000000000000000000000000000000000000000000011110;
  Registers[31] <= 64'b00000000000000000000000000000000000000000000000000000000011111;
  end
  
  always @ (*)
  begin
    if (clk & RegWrite)
      Registers[RD] = WriteData;
    if (reset)
    begin 
      ReadData1 <= 64'b0;
      ReadData2 <= 64'b0;
    end
    else
    begin
      ReadData1 <= Registers[RS1];
      ReadData2 <= Registers[RS2];
    end 
  end
  
endmodule

  
  